module Timeline(
    input [9:0] time_counter,
    output reg [3:0] now
);

    always@(*) begin
        case(time_counter)
            10'd0: now = 4'd8;        10'd1: now = 4'd8;
            10'd2: now = 4'd8;        10'd3: now = 4'd8;
            10'd4: now = 4'd8;        10'd5: now = 4'd1;
            10'd6: now = 4'd1;        10'd7: now = 4'd1;
            10'd8: now = 4'd1;        10'd9: now = 4'd1;
            10'd10: now = 4'd1;        10'd11: now = 4'd1;
            10'd12: now = 4'd1;        10'd13: now = 4'd1;
            10'd14: now = 4'd1;        10'd15: now = 4'd1;
            10'd16: now = 4'd1;        10'd17: now = 4'd1;
            10'd18: now = 4'd1;        10'd19: now = 4'd1;
            10'd20: now = 4'd1;        10'd21: now = 4'd1;
            10'd22: now = 4'd1;        10'd23: now = 4'd1;
            10'd24: now = 4'd1;        10'd25: now = 4'd1;
            10'd26: now = 4'd1;        10'd27: now = 4'd1;
            10'd28: now = 4'd1;        10'd29: now = 4'd1;
            10'd30: now = 4'd1;        10'd31: now = 4'd1;
            10'd32: now = 4'd1;        10'd33: now = 4'd1;
            10'd34: now = 4'd1;        10'd35: now = 4'd1;
            10'd36: now = 4'd1;        10'd37: now = 4'd1;
            10'd38: now = 4'd1;        10'd39: now = 4'd1;
            10'd40: now = 4'd1;        10'd41: now = 4'd1;
            10'd42: now = 4'd1;        10'd43: now = 4'd1;
            10'd44: now = 4'd1;        10'd45: now = 4'd1;
            10'd46: now = 4'd1;        10'd47: now = 4'd1;
            10'd48: now = 4'd1;        10'd49: now = 4'd1;
            10'd50: now = 4'd1;        10'd51: now = 4'd1;
            10'd52: now = 4'd1;        10'd53: now = 4'd1;
            10'd54: now = 4'd1;        10'd55: now = 4'd2;
            10'd56: now = 4'd3;        10'd57: now = 4'd3;
            10'd58: now = 4'd3;        10'd59: now = 4'd3;
            10'd60: now = 4'd3;        10'd61: now = 4'd3;
            10'd62: now = 4'd3;        10'd63: now = 4'd3;
            10'd64: now = 4'd3;        10'd65: now = 4'd3;
            10'd66: now = 4'd3;        10'd67: now = 4'd3;
            10'd68: now = 4'd3;        10'd69: now = 4'd3;
            10'd70: now = 4'd3;        10'd71: now = 4'd3;
            10'd72: now = 4'd3;        10'd73: now = 4'd3;
            10'd74: now = 4'd3;        10'd75: now = 4'd3;
            10'd76: now = 4'd3;        10'd77: now = 4'd3;
            10'd78: now = 4'd3;        10'd79: now = 4'd3;
            10'd80: now = 4'd3;        10'd81: now = 4'd3;
            10'd82: now = 4'd3;        10'd83: now = 4'd3;
            10'd84: now = 4'd3;        10'd85: now = 4'd3;
            10'd86: now = 4'd3;        10'd87: now = 4'd3;
            10'd88: now = 4'd3;        10'd89: now = 4'd3;
            10'd90: now = 4'd3;        10'd91: now = 4'd3;
            10'd92: now = 4'd3;        10'd93: now = 4'd3;
            10'd94: now = 4'd3;        10'd95: now = 4'd3;
            10'd96: now = 4'd3;        10'd97: now = 4'd3;
            10'd98: now = 4'd3;        10'd99: now = 4'd3;
            10'd100: now = 4'd3;        10'd101: now = 4'd3;
            10'd102: now = 4'd0;        10'd103: now = 4'd0;
            10'd104: now = 4'd0;        10'd105: now = 4'd0;
            10'd106: now = 4'd7;        10'd107: now = 4'd0;
            10'd108: now = 4'd0;        10'd109: now = 4'd0;
            10'd110: now = 4'd7;        10'd111: now = 4'd0;
            10'd112: now = 4'd0;        10'd113: now = 4'd7;
            10'd114: now = 4'd0;        10'd115: now = 4'd0;
            10'd116: now = 4'd7;        10'd117: now = 4'd0;
            10'd118: now = 4'd0;        10'd119: now = 4'd7;
            10'd120: now = 4'd0;        10'd121: now = 4'd0;
            10'd122: now = 4'd0;        10'd123: now = 4'd7;
            10'd124: now = 4'd0;        10'd125: now = 4'd0;
            10'd126: now = 4'd7;        10'd127: now = 4'd0;
            10'd128: now = 4'd0;        10'd129: now = 4'd0;
            10'd130: now = 4'd0;        10'd131: now = 4'd0;
            10'd132: now = 4'd7;        10'd133: now = 4'd0;
            10'd134: now = 4'd0;        10'd135: now = 4'd0;
            10'd136: now = 4'd0;        10'd137: now = 4'd0;
            10'd138: now = 4'd0;        10'd139: now = 4'd7;
            10'd140: now = 4'd0;        10'd141: now = 4'd0;
            10'd142: now = 4'd0;        10'd143: now = 4'd0;
            10'd144: now = 4'd0;        10'd145: now = 4'd0;
            10'd146: now = 4'd0;        10'd147: now = 4'd0;
            10'd148: now = 4'd0;        10'd149: now = 4'd0;
            10'd150: now = 4'd0;        10'd151: now = 4'd0;
            10'd152: now = 4'd0;        10'd153: now = 4'd0;
            10'd154: now = 4'd0;        10'd155: now = 4'd3;
            10'd156: now = 4'd3;        10'd157: now = 4'd3;
            10'd158: now = 4'd3;        10'd159: now = 4'd3;
            10'd160: now = 4'd3;        10'd161: now = 4'd3;
            10'd162: now = 4'd3;        10'd163: now = 4'd3;
            10'd164: now = 4'd3;        10'd165: now = 4'd3;
            10'd166: now = 4'd3;        10'd167: now = 4'd3;
            10'd168: now = 4'd3;        10'd169: now = 4'd3;
            10'd170: now = 4'd3;        10'd171: now = 4'd3;
            10'd172: now = 4'd3;        10'd173: now = 4'd3;
            10'd174: now = 4'd3;        10'd175: now = 4'd3;
            10'd176: now = 4'd3;        10'd177: now = 4'd3;
            10'd178: now = 4'd3;        10'd179: now = 4'd3;
            10'd180: now = 4'd3;        10'd181: now = 4'd3;
            10'd182: now = 4'd3;        10'd183: now = 4'd3;
            10'd184: now = 4'd3;        10'd185: now = 4'd3;
            10'd186: now = 4'd3;        10'd187: now = 4'd3;
            10'd188: now = 4'd3;        10'd189: now = 4'd3;
            10'd190: now = 4'd3;        10'd191: now = 4'd3;
            10'd192: now = 4'd3;        10'd193: now = 4'd3;
            10'd194: now = 4'd3;        10'd195: now = 4'd3;
            10'd196: now = 4'd3;        10'd197: now = 4'd3;
            10'd198: now = 4'd3;        10'd199: now = 4'd3;
            10'd200: now = 4'd3;        10'd201: now = 4'd0;
            10'd202: now = 4'd0;        10'd203: now = 4'd7;
            10'd204: now = 4'd0;        10'd205: now = 4'd0;
            10'd206: now = 4'd0;        10'd207: now = 4'd0;
            10'd208: now = 4'd0;        10'd209: now = 4'd7;
            10'd210: now = 4'd0;        10'd211: now = 4'd0;
            10'd212: now = 4'd0;        10'd213: now = 4'd0;
            10'd214: now = 4'd7;        10'd215: now = 4'd0;
            10'd216: now = 4'd0;        10'd217: now = 4'd0;
            10'd218: now = 4'd0;        10'd219: now = 4'd0;
            10'd220: now = 4'd0;        10'd221: now = 4'd0;
            10'd222: now = 4'd0;        10'd223: now = 4'd7;
            10'd224: now = 4'd0;        10'd225: now = 4'd0;
            10'd226: now = 4'd0;        10'd227: now = 4'd0;
            10'd228: now = 4'd0;        10'd229: now = 4'd0;
            10'd230: now = 4'd0;        10'd231: now = 4'd0;
            10'd232: now = 4'd0;        10'd233: now = 4'd0;
            10'd234: now = 4'd0;        10'd235: now = 4'd0;
            10'd236: now = 4'd0;        10'd237: now = 4'd0;
            10'd238: now = 4'd0;        10'd239: now = 4'd4;
            10'd240: now = 4'd4;        10'd241: now = 4'd4;
            10'd242: now = 4'd4;        10'd243: now = 4'd4;
            10'd244: now = 4'd4;        10'd245: now = 4'd4;
            10'd246: now = 4'd4;        10'd247: now = 4'd4;
            10'd248: now = 4'd4;        10'd249: now = 4'd4;
            10'd250: now = 4'd4;        10'd251: now = 4'd4;
            10'd252: now = 4'd4;        10'd253: now = 4'd4;
            10'd254: now = 4'd4;        10'd255: now = 4'd4;
            10'd256: now = 4'd4;        10'd257: now = 4'd4;
            10'd258: now = 4'd4;        10'd259: now = 4'd4;
            10'd260: now = 4'd4;        10'd261: now = 4'd4;
            10'd262: now = 4'd4;        10'd263: now = 4'd4;
            10'd264: now = 4'd4;        10'd265: now = 4'd4;
            10'd266: now = 4'd4;        10'd267: now = 4'd0;
            10'd268: now = 4'd0;        10'd269: now = 4'd7;
            10'd270: now = 4'd0;        10'd271: now = 4'd0;
            10'd272: now = 4'd7;        10'd273: now = 4'd0;
            10'd274: now = 4'd0;        10'd275: now = 4'd0;
            10'd276: now = 4'd0;        10'd277: now = 4'd0;
            10'd278: now = 4'd0;        10'd279: now = 4'd7;
            10'd280: now = 4'd0;        10'd281: now = 4'd0;
            10'd282: now = 4'd0;        10'd283: now = 4'd0;
            10'd284: now = 4'd0;        10'd285: now = 4'd0;
            10'd286: now = 4'd0;        10'd287: now = 4'd0;
            10'd288: now = 4'd0;        10'd289: now = 4'd0;
            10'd290: now = 4'd0;        10'd291: now = 4'd0;
            10'd292: now = 4'd0;        10'd293: now = 4'd0;
            10'd294: now = 4'd0;        10'd295: now = 4'd4;
            10'd296: now = 4'd4;        10'd297: now = 4'd4;
            10'd298: now = 4'd4;        10'd299: now = 4'd4;
            10'd300: now = 4'd4;        10'd301: now = 4'd4;
            10'd302: now = 4'd4;        10'd303: now = 4'd4;
            10'd304: now = 4'd4;        10'd305: now = 4'd4;
            10'd306: now = 4'd4;        10'd307: now = 4'd4;
            10'd308: now = 4'd4;        10'd309: now = 4'd4;
            10'd310: now = 4'd4;        10'd311: now = 4'd4;
            10'd312: now = 4'd4;        10'd313: now = 4'd4;
            10'd314: now = 4'd4;        10'd315: now = 4'd4;
            10'd316: now = 4'd4;        10'd317: now = 4'd4;
            10'd318: now = 4'd4;        10'd319: now = 4'd4;
            10'd320: now = 4'd4;        10'd321: now = 4'd4;
            10'd322: now = 4'd4;        10'd323: now = 4'd0;
            10'd324: now = 4'd0;        10'd325: now = 4'd0;
            10'd326: now = 4'd0;        10'd327: now = 4'd7;
            10'd328: now = 4'd0;        10'd329: now = 4'd0;
            10'd330: now = 4'd0;        10'd331: now = 4'd0;
            10'd332: now = 4'd0;        10'd333: now = 4'd0;
            10'd334: now = 4'd0;        10'd335: now = 4'd0;
            10'd336: now = 4'd0;        10'd337: now = 4'd0;
            10'd338: now = 4'd0;        10'd339: now = 4'd0;
            10'd340: now = 4'd0;        10'd341: now = 4'd0;
            10'd342: now = 4'd0;        10'd343: now = 4'd4;
            10'd344: now = 4'd4;        10'd345: now = 4'd4;
            10'd346: now = 4'd4;        10'd347: now = 4'd4;
            10'd348: now = 4'd4;        10'd349: now = 4'd4;
            10'd350: now = 4'd4;        10'd351: now = 4'd4;
            10'd352: now = 4'd4;        10'd353: now = 4'd4;
            10'd354: now = 4'd4;        10'd355: now = 4'd4;
            10'd356: now = 4'd4;        10'd357: now = 4'd4;
            10'd358: now = 4'd4;        10'd359: now = 4'd4;
            10'd360: now = 4'd4;        10'd361: now = 4'd4;
            10'd362: now = 4'd4;        10'd363: now = 4'd4;
            10'd364: now = 4'd4;        10'd365: now = 4'd4;
            10'd366: now = 4'd4;        10'd367: now = 4'd4;
            10'd368: now = 4'd4;        10'd369: now = 4'd4;
            10'd370: now = 4'd4;        10'd371: now = 4'd0;
            10'd372: now = 4'd0;        10'd373: now = 4'd0;
            10'd374: now = 4'd0;        10'd375: now = 4'd0;
            10'd376: now = 4'd0;        10'd377: now = 4'd0;
            10'd378: now = 4'd0;        10'd379: now = 4'd0;
            10'd380: now = 4'd0;        10'd381: now = 4'd0;
            10'd382: now = 4'd0;        10'd383: now = 4'd0;
            10'd384: now = 4'd0;        10'd385: now = 4'd0;
            10'd386: now = 4'd0;        10'd387: now = 4'd0;
            10'd388: now = 4'd0;        10'd389: now = 4'd0;
            10'd390: now = 4'd0;        10'd391: now = 4'd5;
            10'd392: now = 4'd5;        10'd393: now = 4'd5;
            10'd394: now = 4'd5;        10'd395: now = 4'd5;
            10'd396: now = 4'd5;        10'd397: now = 4'd5;
            10'd398: now = 4'd5;        10'd399: now = 4'd5;
            10'd400: now = 4'd5;        10'd401: now = 4'd5;
            10'd402: now = 4'd5;        10'd403: now = 4'd5;
            10'd404: now = 4'd5;        10'd405: now = 4'd5;
            10'd406: now = 4'd5;        10'd407: now = 4'd5;
            10'd408: now = 4'd5;        10'd409: now = 4'd5;
            10'd410: now = 4'd0;        10'd411: now = 4'd0;
            10'd412: now = 4'd7;        10'd413: now = 4'd0;
            10'd414: now = 4'd0;        10'd415: now = 4'd0;
            10'd416: now = 4'd0;        10'd417: now = 4'd0;
            10'd418: now = 4'd0;        10'd419: now = 4'd0;
            10'd420: now = 4'd0;        10'd421: now = 4'd7;
            10'd422: now = 4'd0;        10'd423: now = 4'd0;
            10'd424: now = 4'd0;        10'd425: now = 4'd0;
            10'd426: now = 4'd0;        10'd427: now = 4'd7;
            10'd428: now = 4'd0;        10'd429: now = 4'd0;
            10'd430: now = 4'd0;        10'd431: now = 4'd0;
            10'd432: now = 4'd0;        10'd433: now = 4'd0;
            10'd434: now = 4'd0;        10'd435: now = 4'd0;
            10'd436: now = 4'd0;        10'd437: now = 4'd0;
            10'd438: now = 4'd0;        10'd439: now = 4'd0;
            10'd440: now = 4'd0;        10'd441: now = 4'd0;
            10'd442: now = 4'd0;        10'd443: now = 4'd5;
            10'd444: now = 4'd5;        10'd445: now = 4'd5;
            10'd446: now = 4'd5;        10'd447: now = 4'd5;
            10'd448: now = 4'd5;        10'd449: now = 4'd5;
            10'd450: now = 4'd5;        10'd451: now = 4'd5;
            10'd452: now = 4'd5;        10'd453: now = 4'd5;
            10'd454: now = 4'd5;        10'd455: now = 4'd5;
            10'd456: now = 4'd5;        10'd457: now = 4'd5;
            10'd458: now = 4'd5;        10'd459: now = 4'd5;
            10'd460: now = 4'd5;        10'd461: now = 4'd5;
            10'd462: now = 4'd0;        10'd463: now = 4'd0;
            10'd464: now = 4'd7;        10'd465: now = 4'd0;
            10'd466: now = 4'd0;        10'd467: now = 4'd0;
            10'd468: now = 4'd0;        10'd469: now = 4'd0;
            10'd470: now = 4'd0;        10'd471: now = 4'd0;
            10'd472: now = 4'd0;        10'd473: now = 4'd0;
            10'd474: now = 4'd0;        10'd475: now = 4'd0;
            10'd476: now = 4'd0;        10'd477: now = 4'd0;
            10'd478: now = 4'd0;        10'd479: now = 4'd0;
            10'd480: now = 4'd6;        10'd481: now = 4'd6;
            10'd482: now = 4'd6;        10'd483: now = 4'd6;
            10'd484: now = 4'd6;        10'd485: now = 4'd6;
            10'd486: now = 4'd6;        10'd487: now = 4'd6;
            10'd488: now = 4'd6;        10'd489: now = 4'd6;
            10'd490: now = 4'd6;        10'd491: now = 4'd6;
            10'd492: now = 4'd0;        10'd493: now = 4'd0;
            10'd494: now = 4'd7;        10'd495: now = 4'd0;
            10'd496: now = 4'd0;        10'd497: now = 4'd7;
            10'd498: now = 4'd0;        10'd499: now = 4'd0;
            10'd500: now = 4'd0;        10'd501: now = 4'd0;
            10'd502: now = 4'd0;        10'd503: now = 4'd7;
            10'd504: now = 4'd0;        10'd505: now = 4'd0;
            10'd506: now = 4'd0;        10'd507: now = 4'd0;
            10'd508: now = 4'd0;        10'd509: now = 4'd0;
            10'd510: now = 4'd7;        10'd511: now = 4'd0;
            10'd512: now = 4'd0;        10'd513: now = 4'd0;
            10'd514: now = 4'd0;        10'd515: now = 4'd0;
            10'd516: now = 4'd0;        10'd517: now = 4'd0;
            10'd518: now = 4'd0;        10'd519: now = 4'd0;
            10'd520: now = 4'd0;        10'd521: now = 4'd0;
            10'd522: now = 4'd0;        10'd523: now = 4'd0;
            10'd524: now = 4'd0;        10'd525: now = 4'd0;
            10'd526: now = 4'd6;        10'd527: now = 4'd6;
            10'd528: now = 4'd6;        10'd529: now = 4'd6;
            10'd530: now = 4'd6;        10'd531: now = 4'd6;
            10'd532: now = 4'd6;        10'd533: now = 4'd6;
            10'd534: now = 4'd6;        10'd535: now = 4'd6;
            10'd536: now = 4'd6;        10'd537: now = 4'd6;
            10'd538: now = 4'd0;        10'd539: now = 4'd0;
            10'd540: now = 4'd0;        10'd541: now = 4'd7;
            10'd542: now = 4'd0;        10'd543: now = 4'd0;
            10'd544: now = 4'd7;        10'd545: now = 4'd0;
            10'd546: now = 4'd0;        10'd547: now = 4'd0;
            10'd548: now = 4'd0;        10'd549: now = 4'd0;
            10'd550: now = 4'd7;        10'd551: now = 4'd0;
            10'd552: now = 4'd0;        10'd553: now = 4'd0;
            10'd554: now = 4'd0;        10'd555: now = 4'd0;
            10'd556: now = 4'd0;        10'd557: now = 4'd0;
            10'd558: now = 4'd0;        10'd559: now = 4'd0;
            10'd560: now = 4'd0;        10'd561: now = 4'd0;
            10'd562: now = 4'd0;        10'd563: now = 4'd0;
            10'd564: now = 4'd0;        10'd565: now = 4'd0;
            10'd566: now = 4'd0;        10'd567: now = 4'd0;
            10'd568: now = 4'd0;        10'd569: now = 4'd0;
            10'd570: now = 4'd0;        10'd571: now = 4'd6;
            10'd572: now = 4'd6;        10'd573: now = 4'd6;
            10'd574: now = 4'd6;        10'd575: now = 4'd6;
            10'd576: now = 4'd6;        10'd577: now = 4'd6;
            10'd578: now = 4'd6;        10'd579: now = 4'd6;
            10'd580: now = 4'd6;        10'd581: now = 4'd6;
            10'd582: now = 4'd6;        default: now = 4'd0;
        endcase
    end

endmodule